type rom_type is array (0 TO 28160) of signed (7 DOWNTO 0);
signal rom : rom_type := (to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), 
to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(37, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(4, 8), to_signed(1, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(41, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(41, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(0, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(0, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(37, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8));