LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY rom_life IS
    PORT (
        CLOCK          : IN  STD_LOGIC;
        ADDR_R         : IN  STD_LOGIC_VECTOR(17 DOWNTO 0);
        DATA_OUT       : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END rom_life;

ARCHITECTURE Behavioral OF rom_life IS
    type rom_type is array (0 TO 2394) of signed (7 DOWNTO 0);
    signal rom : rom_type := (to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(146, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(146, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(0, 8), to_signed(146, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(146, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8),
                              to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8),
                              to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8),
                              to_signed(28, 8), to_signed(28, 8), to_signed(0, 8));
    -- QUELQUES PETITES MODIFICATIONS FAITES POUR AIDER VIVADO A FAIRE LES BONS
    -- CHOIX D'IMPLEMENTATION...

    ATTRIBUTE RAM_STYLE : string;
    ATTRIBUTE RAM_STYLE of rom: signal is "BLOCK";

BEGIN

    PROCESS (CLOCK)
    BEGIN
        IF (CLOCK'event AND CLOCK = '1') THEN
            if unsigned(addr_r) < to_unsigned(2394, 18) then
                DATA_OUT <= STD_LOGIC_VECTOR( rom(to_integer(UNSIGNED(ADDR_R))) );
            end if;
        END IF;
    END PROCESS;

END Behavioral;