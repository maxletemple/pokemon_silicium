type rom_type is array (0 TO 28160) of signed (7 DOWNTO 0);
signal rom : rom_type := (to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), to_signed(122, 8), 
to_signed(122, 8), to_signed(122, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(150, 8), to_signed(150, 8), to_signed(118, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(150, 8), to_signed(150, 8), to_signed(182, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(145, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(109, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(109, 8), to_signed(145, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(145, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(109, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(109, 8), to_signed(145, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(109, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(109, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(109, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(109, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(145, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(109, 8), to_signed(145, 8), to_signed(109, 8), to_signed(109, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(146, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(214, 8), to_signed(218, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(141, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(141, 8), 
to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), 
to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(141, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(178, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(141, 8), to_signed(178, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), to_signed(178, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(178, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(182, 8), to_signed(146, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(178, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(178, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), to_signed(141, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), 
to_signed(214, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(141, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(141, 8), to_signed(178, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(141, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(141, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(141, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(141, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(141, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(141, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(141, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(141, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), 
to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(178, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(178, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(178, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(178, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(178, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(141, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(141, 8), to_signed(69, 8), to_signed(69, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(0, 8));