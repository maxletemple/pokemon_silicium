type rom_type is array (0 TO 8192) of signed (7 DOWNTO 0);
signal rom : rom_type := (to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(46, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), to_signed(82, 8), to_signed(46, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(46, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(82, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), to_signed(82, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(77, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(82, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(255, 8), to_signed(0, 8), to_signed(77, 8), to_signed(255, 8), 
to_signed(82, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(255, 8), to_signed(0, 8), to_signed(0, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(77, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), 
to_signed(255, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(77, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(0, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(77, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(77, 8), to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(0, 8), to_signed(0, 8), to_signed(77, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(77, 8), to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(77, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(140, 8), to_signed(72, 8), to_signed(72, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(77, 8), to_signed(140, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(82, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(46, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), to_signed(9, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(9, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(212, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(136, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(136, 8), to_signed(208, 8), to_signed(249, 8), to_signed(249, 8), 
to_signed(249, 8), to_signed(216, 8), to_signed(216, 8), to_signed(208, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(208, 8), to_signed(249, 8), to_signed(249, 8), to_signed(249, 8), to_signed(249, 8), 
to_signed(249, 8), to_signed(249, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(68, 8), to_signed(208, 8), to_signed(216, 8), to_signed(249, 8), to_signed(249, 8), to_signed(249, 8), to_signed(249, 8), to_signed(249, 8), 
to_signed(249, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(208, 8), 
to_signed(136, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(208, 8), to_signed(0, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(73, 8), to_signed(255, 8), to_signed(0, 8), to_signed(36, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(0, 8), to_signed(255, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(36, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), to_signed(68, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(208, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), 
to_signed(36, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(200, 8), to_signed(200, 8), to_signed(216, 8), 
to_signed(208, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(68, 8), to_signed(136, 8), to_signed(208, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(160, 8), 
to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(200, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(208, 8), to_signed(68, 8), to_signed(136, 8), to_signed(160, 8), to_signed(160, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(208, 8), to_signed(216, 8), to_signed(212, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), 
to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(160, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), 
to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), 
to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(160, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(200, 8), to_signed(200, 8), 
to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(160, 8), to_signed(160, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(200, 8), to_signed(200, 8), 
to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(208, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(208, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(68, 8), to_signed(208, 8), to_signed(208, 8), to_signed(208, 8), 
to_signed(212, 8), to_signed(208, 8), to_signed(68, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(208, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(0, 8), to_signed(208, 8), to_signed(208, 8), to_signed(208, 8), to_signed(208, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(208, 8), to_signed(208, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(0, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(208, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(0, 8), to_signed(216, 8), to_signed(208, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(68, 8), to_signed(136, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(216, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(208, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(208, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(68, 8), to_signed(136, 8), to_signed(136, 8), to_signed(208, 8), 
to_signed(208, 8), to_signed(136, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(216, 8), to_signed(136, 8), 
to_signed(216, 8), to_signed(208, 8), to_signed(68, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8));