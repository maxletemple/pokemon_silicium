type rom_type IS array (0 TO 9497) OF SIGNED (7 DOWNTO 0);
signal rom : rom_type := (to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(217, 8), to_signed(73, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(172, 8), to_signed(217, 8), to_signed(217, 8), to_signed(216, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(172, 8), to_signed(217, 8), to_signed(217, 8), to_signed(216, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(212, 8), to_signed(172, 8), 
to_signed(172, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(104, 8), to_signed(0, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(172, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(172, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(212, 8), to_signed(172, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(212, 8), 
to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(0, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), 
to_signed(172, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(104, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(104, 8), to_signed(104, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(172, 8), to_signed(217, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), 
to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(172, 8), to_signed(104, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(46, 8), to_signed(104, 8), to_signed(217, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), 
to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(216, 8), to_signed(172, 8), to_signed(172, 8), to_signed(216, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(216, 8), to_signed(217, 8), 
to_signed(216, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(104, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(216, 8), to_signed(217, 8), to_signed(216, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(172, 8), to_signed(212, 8), to_signed(212, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(217, 8), to_signed(216, 8), to_signed(217, 8), 
to_signed(216, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(104, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(172, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(172, 8), to_signed(172, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(217, 8), to_signed(216, 8), to_signed(217, 8), to_signed(216, 8), to_signed(217, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(172, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(212, 8), to_signed(217, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(172, 8), to_signed(172, 8), to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(172, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(212, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(172, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(104, 8), 
to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(104, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(212, 8), to_signed(196, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(172, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(192, 8), to_signed(196, 8), to_signed(0, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(172, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), 
to_signed(192, 8), to_signed(192, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(104, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(192, 8), to_signed(192, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(217, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(172, 8), to_signed(192, 8), 
to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(104, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(172, 8), to_signed(104, 8), to_signed(172, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(172, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(104, 8), to_signed(104, 8), to_signed(216, 8), to_signed(172, 8), to_signed(172, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(217, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(172, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(172, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(172, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(217, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(0, 8), to_signed(172, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(172, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(104, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(217, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(104, 8), 
to_signed(172, 8), to_signed(104, 8), to_signed(172, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(172, 8), to_signed(172, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(104, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(217, 8), to_signed(216, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(172, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(104, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(104, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(104, 8), to_signed(212, 8), to_signed(172, 8), to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(216, 8), to_signed(0, 8), to_signed(172, 8), to_signed(172, 8), 
to_signed(172, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(172, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(172, 8), 
to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(172, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(172, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(104, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(9, 8), to_signed(82, 8), to_signed(46, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(82, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(82, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), to_signed(82, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(255, 8), to_signed(255, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(255, 8), to_signed(0, 8), to_signed(0, 8), to_signed(255, 8), 
to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), 
to_signed(77, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), 
to_signed(77, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(0, 8), to_signed(182, 8), to_signed(77, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(0, 8), to_signed(0, 8), to_signed(77, 8), to_signed(182, 8), 
to_signed(77, 8), to_signed(212, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(182, 8), to_signed(182, 8), to_signed(72, 8), to_signed(72, 8), to_signed(0, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(140, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(46, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), 
to_signed(82, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(0, 8), to_signed(9, 8), to_signed(46, 8), to_signed(0, 8), to_signed(46, 8), to_signed(0, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(46, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(150, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(9, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(46, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), 
to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), to_signed(101, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), to_signed(101, 8), to_signed(137, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), to_signed(174, 8), 
to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(101, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), to_signed(101, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(137, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(36, 8), to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), 
to_signed(101, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(101, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(137, 8), to_signed(36, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), 
to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(36, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), to_signed(174, 8), to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(36, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), to_signed(101, 8), to_signed(137, 8), 
to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(101, 8), to_signed(36, 8), to_signed(36, 8), to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(137, 8), to_signed(0, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(36, 8), to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(0, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(36, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), 
to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(0, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(0, 8), to_signed(101, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(137, 8), 
to_signed(137, 8), to_signed(101, 8), to_signed(36, 8), to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), to_signed(0, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), 
to_signed(101, 8), to_signed(36, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(0, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(101, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(164, 8), to_signed(36, 8), to_signed(101, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), 
to_signed(174, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(200, 8), to_signed(164, 8), to_signed(36, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(200, 8), to_signed(209, 8), to_signed(164, 8), 
to_signed(101, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), 
to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(200, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(200, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(200, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(36, 8), to_signed(101, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(200, 8), to_signed(200, 8), 
to_signed(36, 8), to_signed(101, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(0, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(200, 8), to_signed(200, 8), 
to_signed(200, 8), to_signed(101, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), 
to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(182, 8), to_signed(174, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(200, 8), 
to_signed(200, 8), to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(0, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(36, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(182, 8), to_signed(182, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(36, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(174, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(174, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(101, 8), to_signed(174, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(174, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(101, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(109, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(109, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(36, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(218, 8), to_signed(218, 8), to_signed(109, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(109, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(36, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(218, 8), to_signed(218, 8), to_signed(109, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(218, 8), to_signed(109, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(36, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(109, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), to_signed(36, 8), to_signed(36, 8), to_signed(101, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(101, 8), to_signed(36, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(36, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(109, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(36, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(0, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), 
to_signed(36, 8), to_signed(101, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(137, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(137, 8), to_signed(36, 8), to_signed(36, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(137, 8), to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(137, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(36, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(137, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(137, 8), to_signed(137, 8), to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(0, 8));