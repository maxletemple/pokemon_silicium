type rom_type is array(0 to 577) of unsigned(6 downto 0); 
 signal rom : rom_type := (to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(4, 7),to_unsigned(28, 7),to_unsigned(45, 7),to_unsigned(40, 7),to_unsigned(41, 7),to_unsigned(37, 7),to_unsigned(26, 7),to_unsigned(44, 7),to_unsigned(38, 7),to_unsigned(26, 7),
to_unsigned(19, 7),to_unsigned(34, 7),to_unsigned(41, 7),to_unsigned(37, 7),to_unsigned(40, 7),to_unsigned(46, 7),to_unsigned(31, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(15, 7),to_unsigned(34, 7),to_unsigned(36, 7),to_unsigned(26, 7),to_unsigned(28, 7),to_unsigned(33, 7),to_unsigned(46, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(1, 7),to_unsigned(43, 7),to_unsigned(26, 7),to_unsigned(44, 7),to_unsigned(66, 7), to_unsigned(32, 7),to_unsigned(26, 7),to_unsigned(37, 7),to_unsigned(34, 7),to_unsigned(69, 7), 
to_unsigned(19, 7),to_unsigned(40, 7),to_unsigned(43, 7),to_unsigned(45, 7),to_unsigned(30, 7),to_unsigned(43, 7),to_unsigned(43, 7),to_unsigned(26, 7),to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(17, 7),to_unsigned(26, 7),to_unsigned(50, 7),to_unsigned(42, 7),to_unsigned(46, 7),to_unsigned(26, 7),to_unsigned(51, 7),to_unsigned(26, 7),to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(12, 7),to_unsigned(30, 7),to_unsigned(48, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(17, 7),to_unsigned(40, 7),to_unsigned(39, 7),to_unsigned(31, 7),to_unsigned(37, 7),to_unsigned(30, 7),to_unsigned(49, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(1, 7),to_unsigned(40, 7),to_unsigned(38, 7),to_unsigned(27, 7),to_unsigned(43, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(6, 7),to_unsigned(26, 7),to_unsigned(51, 7),to_unsigned(69, 7), to_unsigned(19, 7),to_unsigned(40, 7),to_unsigned(49, 7),to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(11, 7),to_unsigned(26, 7),to_unsigned(43, 7),to_unsigned(28, 7),to_unsigned(34, 7),to_unsigned(39, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(8, 7),to_unsigned(38, 7),to_unsigned(41, 7),to_unsigned(26, 7),to_unsigned(28, 7),to_unsigned(45, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(15, 7),to_unsigned(34, 7),to_unsigned(28, 7),to_unsigned(26, 7),to_unsigned(43, 7),to_unsigned(29, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(15, 7),to_unsigned(34, 7),to_unsigned(28, 7),to_unsigned(41, 7),to_unsigned(34, 7),to_unsigned(28, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(2, 7),to_unsigned(33, 7),to_unsigned(26, 7),to_unsigned(43, 7),to_unsigned(32, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(18, 7),to_unsigned(46, 7),to_unsigned(43, 7),to_unsigned(31, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(4, 7),to_unsigned(28, 7),to_unsigned(37, 7),to_unsigned(26, 7),to_unsigned(34, 7),to_unsigned(43, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(10, 7),to_unsigned(30, 7),to_unsigned(46, 7),to_unsigned(29, 7),to_unsigned(31, 7),to_unsigned(30, 7),to_unsigned(43, 7),to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(4, 7),to_unsigned(28, 7),to_unsigned(37, 7),to_unsigned(26, 7),to_unsigned(45, 7),to_unsigned(43, 7),to_unsigned(40, 7),to_unsigned(28, 7),to_unsigned(69, 7), 
to_unsigned(19, 7),to_unsigned(46, 7),to_unsigned(39, 7),to_unsigned(39, 7),to_unsigned(30, 7),to_unsigned(37, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(6, 7),to_unsigned(43, 7),to_unsigned(34, 7),to_unsigned(31, 7),to_unsigned(31, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(7, 7),to_unsigned(34, 7),to_unsigned(32, 7),to_unsigned(33, 7),to_unsigned(69, 7), to_unsigned(10, 7),to_unsigned(34, 7),to_unsigned(36, 7),to_unsigned(69, 7), 
to_unsigned(12, 7),to_unsigned(40, 7),to_unsigned(37, 7),to_unsigned(40, 7),to_unsigned(45, 7),to_unsigned(40, 7),to_unsigned(47, 7),to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(21, 7),to_unsigned(30, 7),to_unsigned(39, 7),to_unsigned(29, 7),to_unsigned(30, 7),to_unsigned(45, 7),to_unsigned(45, 7),to_unsigned(26, 7),to_unsigned(69, 7), 
to_unsigned(18, 7),to_unsigned(66, 7), to_unsigned(34, 7),to_unsigned(44, 7),to_unsigned(38, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(2, 7),to_unsigned(33, 7),to_unsigned(26, 7),to_unsigned(39, 7),to_unsigned(47, 7),to_unsigned(43, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(12, 7),to_unsigned(40, 7),to_unsigned(43, 7),to_unsigned(44, 7),to_unsigned(46, 7),to_unsigned(43, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(19, 7),to_unsigned(26, 7),to_unsigned(41, 7),to_unsigned(40, 7),to_unsigned(45, 7),to_unsigned(34, 7),to_unsigned(32, 7),to_unsigned(30, 7),to_unsigned(69, 7), 
to_unsigned(14, 7),to_unsigned(46, 7),to_unsigned(43, 7),to_unsigned(26, 7),to_unsigned(32, 7),to_unsigned(26, 7),to_unsigned(39, 7),to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(2, 7),to_unsigned(40, 7),to_unsigned(37, 7),to_unsigned(65, 7), to_unsigned(43, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(3, 7),to_unsigned(43, 7),to_unsigned(26, 7),to_unsigned(28, 7),to_unsigned(40, 7),to_unsigned(43, 7),to_unsigned(26, 7),to_unsigned(32, 7),to_unsigned(30, 7),
to_unsigned(21, 7),to_unsigned(40, 7),to_unsigned(37, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(15, 7),to_unsigned(44, 7),to_unsigned(50, 7),to_unsigned(36, 7),to_unsigned(40, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(4, 7),to_unsigned(39, 7),to_unsigned(45, 7),to_unsigned(43, 7),to_unsigned(26, 7),to_unsigned(47, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(3, 7),to_unsigned(40, 7),to_unsigned(46, 7),to_unsigned(29, 7),to_unsigned(40, 7),to_unsigned(46, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(1, 7),to_unsigned(43, 7),to_unsigned(46, 7),to_unsigned(38, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(2, 7),to_unsigned(33, 7),to_unsigned(26, 7),to_unsigned(43, 7),to_unsigned(32, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(1, 7),to_unsigned(26, 7),to_unsigned(37, 7),to_unsigned(40, 7),to_unsigned(38, 7),to_unsigned(27, 7),to_unsigned(43, 7),to_unsigned(30, 7),to_unsigned(69, 7), 
to_unsigned(6, 7),to_unsigned(34, 7),to_unsigned(31, 7),to_unsigned(37, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(2, 7),to_unsigned(40, 7),to_unsigned(28, 7),to_unsigned(33, 7),to_unsigned(38, 7),to_unsigned(26, 7),to_unsigned(43, 7),to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(0, 7),to_unsigned(45, 7),to_unsigned(45, 7),to_unsigned(26, 7),to_unsigned(42, 7),to_unsigned(46, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(14, 7),to_unsigned(27, 7),to_unsigned(35, 7),to_unsigned(30, 7),to_unsigned(45, 7),to_unsigned(44, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(15, 7),to_unsigned(40, 7),to_unsigned(36, 7),to_unsigned(66, 7), to_unsigned(38, 7),to_unsigned(40, 7),to_unsigned(39, 7),to_unsigned(44, 7),to_unsigned(69, 7), 
to_unsigned(5, 7),to_unsigned(46, 7),to_unsigned(34, 7),to_unsigned(45, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), to_unsigned(69, 7), 
to_unsigned(2, 7),to_unsigned(67, 7), to_unsigned(30, 7),to_unsigned(44, 7),to_unsigned(45, 7),to_unsigned(69, 7), to_unsigned(30, 7),to_unsigned(31, 7),to_unsigned(31, 7),to_unsigned(34, 7),to_unsigned(28, 7),to_unsigned(26, 7),to_unsigned(28, 7),to_unsigned(30, 7),
to_unsigned(2, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(39, 7),to_unsigned(67, 7), to_unsigned(30, 7),to_unsigned(44, 7),to_unsigned(45, 7),to_unsigned(69, 7), to_unsigned(41, 7),to_unsigned(26, 7),to_unsigned(44, 7),to_unsigned(69, 7), to_unsigned(45, 7),to_unsigned(43, 7),to_unsigned(65, 7), to_unsigned(44, 7),to_unsigned(69, 7), to_unsigned(30, 7),to_unsigned(31, 7),to_unsigned(31, 7),to_unsigned(34, 7),to_unsigned(28, 7),to_unsigned(26, 7),to_unsigned(28, 7),to_unsigned(30, 7),
to_unsigned(0, 7),to_unsigned(45, 7),to_unsigned(45, 7),to_unsigned(26, 7),to_unsigned(42, 7),to_unsigned(46, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(28, 7),to_unsigned(40, 7),to_unsigned(43, 7),to_unsigned(43, 7),to_unsigned(30, 7),to_unsigned(28, 7),to_unsigned(45, 7),to_unsigned(30, 7),
to_unsigned(1, 7),to_unsigned(34, 7),to_unsigned(30, 7),to_unsigned(39, 7),to_unsigned(47, 7),to_unsigned(30, 7),to_unsigned(39, 7),to_unsigned(46, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(29, 7),to_unsigned(26, 7),to_unsigned(39, 7),to_unsigned(44, 7),
to_unsigned(41, 7),to_unsigned(40, 7),to_unsigned(36, 7),to_unsigned(66, 7), to_unsigned(38, 7),to_unsigned(40, 7),to_unsigned(39, 7),to_unsigned(69, 7), to_unsigned(44, 7),to_unsigned(34, 7),to_unsigned(37, 7),to_unsigned(34, 7),to_unsigned(28, 7),to_unsigned(34, 7),to_unsigned(46, 7),to_unsigned(38, 7),
to_unsigned(2, 7),to_unsigned(33, 7),to_unsigned(40, 7),to_unsigned(34, 7),to_unsigned(44, 7),to_unsigned(34, 7),to_unsigned(44, 7),to_unsigned(44, 7),to_unsigned(30, 7),to_unsigned(51, 7),
to_unsigned(15, 7),to_unsigned(26, 7),to_unsigned(44, 7),to_unsigned(69, 7), to_unsigned(34, 7),to_unsigned(38, 7),to_unsigned(41, 7),to_unsigned(37, 7),to_unsigned(66, 7), to_unsigned(38, 7),to_unsigned(30, 7),to_unsigned(39, 7),to_unsigned(45, 7),to_unsigned(66, 7), 
to_unsigned(14, 7),to_unsigned(39, 7),to_unsigned(69, 7), to_unsigned(39, 7),to_unsigned(30, 7),to_unsigned(69, 7), to_unsigned(31, 7),to_unsigned(46, 7),to_unsigned(34, 7),to_unsigned(45, 7),to_unsigned(69, 7), to_unsigned(41, 7),to_unsigned(26, 7),to_unsigned(44, 7),
to_unsigned(37, 7),to_unsigned(40, 7),to_unsigned(43, 7),to_unsigned(44, 7),to_unsigned(69, 7), to_unsigned(29, 7),to_unsigned(67, 7), to_unsigned(46, 7),to_unsigned(39, 7),to_unsigned(69, 7), to_unsigned(28, 7),to_unsigned(40, 7),to_unsigned(38, 7),to_unsigned(27, 7),to_unsigned(26, 7),to_unsigned(45, 7),
to_unsigned(0, 7));