type rom_type is array (0 TO 65536) of signed (7 DOWNTO 0);
signal rom : rom_type := (to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(73, 8), to_signed(37, 8), to_signed(37, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(37, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(37, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), 
to_signed(110, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(110, 8), 
to_signed(110, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(37, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(110, 8), to_signed(110, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(37, 8), to_signed(37, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(73, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(110, 8), to_signed(110, 8), to_signed(109, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(73, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(37, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(110, 8), to_signed(110, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(37, 8), to_signed(73, 8), 
to_signed(110, 8), to_signed(110, 8), to_signed(110, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(110, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(109, 8), to_signed(110, 8), to_signed(110, 8), to_signed(110, 8), 
to_signed(110, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(37, 8), to_signed(37, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(217, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(213, 8), to_signed(217, 8), to_signed(144, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(144, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(144, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(144, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(144, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(144, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), 
to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(73, 8), to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(37, 8), to_signed(37, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(37, 8), to_signed(37, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(37, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(110, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(37, 8), to_signed(110, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(110, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(73, 8), to_signed(110, 8), to_signed(110, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(37, 8), to_signed(110, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(37, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(37, 8), to_signed(110, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(113, 8), to_signed(77, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(113, 8), to_signed(113, 8), to_signed(77, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(113, 8), to_signed(113, 8), to_signed(113, 8), 
to_signed(77, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(40, 8), to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(113, 8), 
to_signed(113, 8), to_signed(113, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(40, 8), 
to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(73, 8), to_signed(73, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(113, 8), to_signed(113, 8), to_signed(113, 8), to_signed(77, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(217, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(0, 8), to_signed(0, 8), to_signed(218, 8), 
to_signed(113, 8), to_signed(113, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(0, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(177, 8), to_signed(108, 8), 
to_signed(108, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(108, 8), to_signed(108, 8), to_signed(108, 8), to_signed(177, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(0, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(113, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(177, 8), to_signed(108, 8), to_signed(108, 8), to_signed(217, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), 
to_signed(108, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(113, 8), to_signed(77, 8), 
to_signed(77, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(177, 8), to_signed(108, 8), to_signed(217, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(0, 8), to_signed(108, 8), to_signed(160, 8), to_signed(160, 8), to_signed(218, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(113, 8), to_signed(113, 8), to_signed(77, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(108, 8), to_signed(213, 8), to_signed(217, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(77, 8), to_signed(77, 8), to_signed(113, 8), to_signed(113, 8), to_signed(77, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(108, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(108, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), 
to_signed(160, 8), to_signed(160, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(217, 8), to_signed(113, 8), to_signed(77, 8), to_signed(77, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(108, 8), to_signed(160, 8), to_signed(160, 8), 
to_signed(160, 8), to_signed(160, 8), to_signed(218, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(73, 8), to_signed(217, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(160, 8), 
to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(160, 8), 
to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(77, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), 
to_signed(160, 8), to_signed(160, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(77, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(40, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(77, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(77, 8), to_signed(40, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(77, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(40, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(77, 8), to_signed(40, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(40, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(77, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(0, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(77, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(77, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(73, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(218, 8), to_signed(73, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(77, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(218, 8), to_signed(218, 8), to_signed(108, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(73, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(73, 8), to_signed(218, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), to_signed(218, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(40, 8), to_signed(0, 8), to_signed(218, 8), to_signed(0, 8), to_signed(77, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(77, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(182, 8), to_signed(218, 8), to_signed(0, 8), to_signed(73, 8), to_signed(0, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(0, 8), to_signed(218, 8), to_signed(218, 8), to_signed(0, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(73, 8), to_signed(182, 8), to_signed(73, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(0, 8), to_signed(218, 8), to_signed(182, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(73, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(40, 8), to_signed(218, 8), to_signed(77, 8), 
to_signed(73, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(77, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(77, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(40, 8), to_signed(0, 8), to_signed(40, 8), 
to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(108, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(77, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(40, 8), to_signed(218, 8), to_signed(77, 8), 
to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(73, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(77, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(213, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(213, 8), 
to_signed(73, 8), to_signed(218, 8), to_signed(73, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(77, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(218, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(108, 8), to_signed(213, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(0, 8), to_signed(218, 8), to_signed(0, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(177, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(0, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(0, 8), to_signed(77, 8), to_signed(40, 8), to_signed(40, 8), to_signed(73, 8), 
to_signed(218, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(0, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(77, 8), to_signed(40, 8), to_signed(0, 8), 
to_signed(218, 8), to_signed(182, 8), to_signed(218, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(77, 8), to_signed(0, 8), to_signed(217, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(0, 8), to_signed(213, 8), to_signed(217, 8), to_signed(0, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(177, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(73, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(73, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(108, 8), to_signed(213, 8), to_signed(172, 8), to_signed(172, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(73, 8), 
to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(108, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(73, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(108, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), 
to_signed(172, 8), to_signed(172, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(0, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(172, 8), 
to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(172, 8), to_signed(172, 8), 
to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(172, 8), to_signed(172, 8), 
to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(108, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(108, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(172, 8), 
to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(172, 8), 
to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(172, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(177, 8), to_signed(172, 8), to_signed(172, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(108, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(108, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(108, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(108, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(128, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(164, 8), to_signed(128, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(164, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(164, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(164, 8), to_signed(164, 8), to_signed(128, 8), to_signed(128, 8), to_signed(36, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(164, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(164, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(128, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(164, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(164, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(128, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(128, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(205, 8), to_signed(205, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(205, 8), to_signed(128, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(28, 8), to_signed(128, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(128, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(205, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(205, 8), to_signed(128, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), 
to_signed(128, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), 
to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(128, 8), 
to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(128, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), 
to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(128, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(128, 8), to_signed(205, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(205, 8), to_signed(128, 8), to_signed(128, 8), 
to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(128, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(205, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(36, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(128, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), 
to_signed(128, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(128, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(205, 8), to_signed(128, 8), to_signed(36, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), 
to_signed(214, 8), to_signed(128, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(164, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), 
to_signed(128, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(128, 8), to_signed(36, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(205, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(205, 8), to_signed(128, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(205, 8), to_signed(205, 8), 
to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(128, 8), to_signed(205, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(205, 8), to_signed(128, 8), 
to_signed(128, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(128, 8), to_signed(128, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(128, 8), to_signed(128, 8), to_signed(128, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(128, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), 
to_signed(205, 8), to_signed(128, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(205, 8), to_signed(128, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(205, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(128, 8), to_signed(128, 8), to_signed(205, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(205, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(205, 8), to_signed(164, 8), to_signed(164, 8), to_signed(205, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(214, 8), to_signed(214, 8), to_signed(205, 8), to_signed(164, 8), 
to_signed(164, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(164, 8), to_signed(164, 8), to_signed(164, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(205, 8), to_signed(164, 8), to_signed(164, 8), 
to_signed(164, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(128, 8), to_signed(205, 8), to_signed(164, 8), to_signed(164, 8), to_signed(164, 8), to_signed(205, 8), to_signed(128, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(205, 8), to_signed(164, 8), to_signed(164, 8), 
to_signed(164, 8), to_signed(205, 8), to_signed(128, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(205, 8), to_signed(205, 8), to_signed(164, 8), to_signed(164, 8), to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(205, 8), to_signed(164, 8), 
to_signed(164, 8), to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(128, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(128, 8), to_signed(205, 8), to_signed(205, 8), 
to_signed(205, 8), to_signed(205, 8), to_signed(205, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(164, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(164, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(164, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(164, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(209, 8), to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(164, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(164, 8), to_signed(132, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), to_signed(132, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(164, 8), to_signed(214, 8), to_signed(214, 8), to_signed(132, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(164, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(164, 8), to_signed(214, 8), to_signed(36, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(132, 8), to_signed(173, 8), to_signed(173, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(164, 8), 
to_signed(164, 8), to_signed(209, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(164, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(173, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(164, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(173, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(132, 8), to_signed(164, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(132, 8), to_signed(173, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(132, 8), to_signed(164, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(218, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(36, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(209, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(9, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(164, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(9, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), to_signed(132, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(209, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(36, 8), to_signed(218, 8), to_signed(82, 8), to_signed(218, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(132, 8), to_signed(9, 8), to_signed(82, 8), to_signed(218, 8), to_signed(218, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(132, 8), 
to_signed(214, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(209, 8), to_signed(214, 8), 
to_signed(132, 8), to_signed(9, 8), to_signed(9, 8), to_signed(218, 8), to_signed(218, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(214, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(214, 8), to_signed(164, 8), to_signed(164, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(132, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(132, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(164, 8), to_signed(132, 8), to_signed(132, 8), to_signed(36, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(214, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(173, 8), to_signed(173, 8), to_signed(173, 8), to_signed(173, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(132, 8), to_signed(164, 8), to_signed(164, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(214, 8), 
to_signed(164, 8), to_signed(214, 8), to_signed(214, 8), to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(214, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(132, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(132, 8), to_signed(132, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), 
to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), 
to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(214, 8), to_signed(209, 8), to_signed(164, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(209, 8), to_signed(132, 8), to_signed(209, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(209, 8), to_signed(36, 8), to_signed(132, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(164, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(132, 8), 
to_signed(209, 8), to_signed(36, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(214, 8), to_signed(209, 8), 
to_signed(164, 8), to_signed(36, 8), to_signed(214, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(164, 8), to_signed(132, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(132, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(164, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(214, 8), to_signed(164, 8), 
to_signed(164, 8), to_signed(36, 8), to_signed(214, 8), to_signed(132, 8), to_signed(209, 8), to_signed(209, 8), to_signed(164, 8), to_signed(36, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(214, 8), 
to_signed(209, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(164, 8), 
to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(132, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(214, 8), to_signed(209, 8), to_signed(164, 8), 
to_signed(36, 8), to_signed(173, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(164, 8), to_signed(209, 8), to_signed(214, 8), to_signed(214, 8), to_signed(132, 8), to_signed(214, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(36, 8), to_signed(173, 8), to_signed(132, 8), to_signed(132, 8), to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(132, 8), 
to_signed(173, 8), to_signed(173, 8), to_signed(36, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(132, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), 
to_signed(173, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(132, 8), to_signed(214, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(173, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(132, 8), to_signed(209, 8), to_signed(173, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), 
to_signed(214, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(132, 8), to_signed(173, 8), to_signed(173, 8), to_signed(173, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(173, 8), 
to_signed(173, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(132, 8), to_signed(214, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(173, 8), to_signed(173, 8), to_signed(132, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(209, 8), to_signed(209, 8), to_signed(132, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(132, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(132, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(214, 8), to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(132, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(45, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(45, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(118, 8), 
to_signed(85, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(45, 8), to_signed(85, 8), to_signed(118, 8), to_signed(85, 8), 
to_signed(118, 8), to_signed(85, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(0, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(118, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(180, 8), to_signed(216, 8), to_signed(180, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(118, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(180, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), 
to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(216, 8), to_signed(216, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(118, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(216, 8), to_signed(216, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(173, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(216, 8), to_signed(180, 8), to_signed(118, 8), to_signed(180, 8), to_signed(180, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(173, 8), to_signed(201, 8), to_signed(201, 8), to_signed(173, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(216, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(216, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(173, 8), to_signed(201, 8), to_signed(201, 8), to_signed(201, 8), to_signed(201, 8), to_signed(173, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(180, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(85, 8), to_signed(118, 8), to_signed(85, 8), to_signed(118, 8), to_signed(180, 8), to_signed(180, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(201, 8), to_signed(201, 8), to_signed(45, 8), to_signed(40, 8), to_signed(201, 8), to_signed(201, 8), 
to_signed(201, 8), to_signed(85, 8), to_signed(40, 8), to_signed(216, 8), to_signed(0, 8), to_signed(118, 8), to_signed(45, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(45, 8), to_signed(118, 8), to_signed(85, 8), 
to_signed(118, 8), to_signed(85, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(201, 8), to_signed(40, 8), to_signed(41, 8), to_signed(41, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(201, 8), to_signed(201, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(201, 8), to_signed(40, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(201, 8), to_signed(173, 8), to_signed(85, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(85, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(173, 8), to_signed(201, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(40, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(40, 8), to_signed(40, 8), to_signed(173, 8), to_signed(118, 8), to_signed(118, 8), to_signed(45, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(173, 8), to_signed(201, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(40, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(173, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(41, 8), to_signed(41, 8), to_signed(40, 8), to_signed(40, 8), to_signed(118, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(180, 8), to_signed(180, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(173, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(182, 8), to_signed(40, 8), to_signed(41, 8), to_signed(40, 8), to_signed(85, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(45, 8), to_signed(173, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(28, 8), to_signed(40, 8), to_signed(218, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(180, 8), to_signed(180, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(173, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(173, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(180, 8), to_signed(180, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(173, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(45, 8), to_signed(173, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(173, 8), to_signed(173, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(45, 8), to_signed(173, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(180, 8), to_signed(180, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(180, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(180, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(180, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(180, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(0, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(218, 8), to_signed(218, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(182, 8), to_signed(182, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(218, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(45, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(182, 8), to_signed(182, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(85, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(40, 8), to_signed(118, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(216, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(118, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(180, 8), to_signed(180, 8), to_signed(40, 8), to_signed(118, 8), 
to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(118, 8), to_signed(85, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(40, 8), to_signed(118, 8), to_signed(85, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(44, 8), to_signed(44, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), 
to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(180, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(44, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(201, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(44, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(180, 8), to_signed(180, 8), to_signed(40, 8), to_signed(40, 8), to_signed(44, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(216, 8), 
to_signed(180, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(201, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(44, 8), to_signed(44, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(44, 8), to_signed(0, 8), to_signed(216, 8), to_signed(40, 8), to_signed(44, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(216, 8), to_signed(180, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(201, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(44, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(173, 8), to_signed(201, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(216, 8), to_signed(180, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(201, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(173, 8), to_signed(173, 8), to_signed(173, 8), to_signed(173, 8), to_signed(173, 8), to_signed(173, 8), to_signed(173, 8), 
to_signed(173, 8), to_signed(201, 8), to_signed(201, 8), to_signed(201, 8), to_signed(201, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(180, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(201, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(218, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(201, 8), to_signed(201, 8), to_signed(173, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(180, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(85, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(201, 8), to_signed(201, 8), to_signed(201, 8), to_signed(201, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(40, 8), to_signed(201, 8), to_signed(173, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(180, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(118, 8), to_signed(45, 8), to_signed(40, 8), to_signed(201, 8), 
to_signed(201, 8), to_signed(201, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(0, 8), to_signed(201, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), 
to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(180, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(0, 8), to_signed(201, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(0, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(0, 8), to_signed(201, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(50, 8), 
to_signed(41, 8), to_signed(40, 8), to_signed(201, 8), to_signed(173, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(0, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(85, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(50, 8), to_signed(50, 8), 
to_signed(50, 8), to_signed(0, 8), to_signed(201, 8), to_signed(45, 8), to_signed(0, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(45, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(45, 8), to_signed(85, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(50, 8), to_signed(50, 8), to_signed(50, 8), 
to_signed(40, 8), to_signed(201, 8), to_signed(173, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(45, 8), 
to_signed(85, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(50, 8), to_signed(50, 8), to_signed(41, 8), 
to_signed(0, 8), to_signed(173, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(85, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), 
to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(173, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(173, 8), to_signed(45, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(0, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(40, 8), to_signed(85, 8), to_signed(40, 8), to_signed(85, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(173, 8), to_signed(173, 8), to_signed(173, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), 
to_signed(40, 8), to_signed(218, 8), to_signed(218, 8), to_signed(45, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(0, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(0, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(0, 8), to_signed(85, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(40, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(45, 8), to_signed(85, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(0, 8), to_signed(85, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(0, 8), to_signed(40, 8), to_signed(182, 8), 
to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(218, 8), to_signed(218, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(40, 8), 
to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(45, 8), to_signed(0, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(40, 8), to_signed(201, 8), to_signed(201, 8), to_signed(40, 8), to_signed(218, 8), to_signed(0, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(85, 8), to_signed(40, 8), to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), 
to_signed(0, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), to_signed(0, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(45, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(218, 8), to_signed(218, 8), to_signed(0, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(0, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(40, 8), to_signed(40, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(40, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), 
to_signed(0, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(173, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(0, 8), to_signed(28, 8), to_signed(40, 8), to_signed(0, 8), to_signed(182, 8), to_signed(0, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(85, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(173, 8), to_signed(0, 8), to_signed(0, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(44, 8), to_signed(0, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(173, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(0, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(201, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(0, 8), to_signed(45, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(201, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(45, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(201, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), to_signed(118, 8), to_signed(85, 8), to_signed(118, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(201, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(180, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(180, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), to_signed(85, 8), to_signed(118, 8), to_signed(85, 8), 
to_signed(118, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(201, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(180, 8), to_signed(216, 8), to_signed(180, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(180, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), to_signed(85, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(201, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(180, 8), to_signed(45, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(40, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(180, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), 
to_signed(201, 8), to_signed(201, 8), to_signed(201, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(216, 8), to_signed(180, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(201, 8), to_signed(201, 8), to_signed(201, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), 
to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(216, 8), to_signed(180, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(40, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(201, 8), to_signed(201, 8), 
to_signed(201, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(118, 8), to_signed(118, 8), to_signed(45, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(180, 8), to_signed(216, 8), to_signed(216, 8), to_signed(85, 8), to_signed(216, 8), 
to_signed(180, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(201, 8), to_signed(201, 8), to_signed(201, 8), to_signed(118, 8), to_signed(118, 8), to_signed(85, 8), to_signed(201, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(118, 8), to_signed(40, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(40, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(201, 8), to_signed(201, 8), to_signed(201, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(118, 8), to_signed(40, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(85, 8), 
to_signed(85, 8), to_signed(216, 8), to_signed(85, 8), to_signed(85, 8), to_signed(216, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(40, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(85, 8), to_signed(201, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(173, 8), to_signed(85, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(118, 8), to_signed(45, 8), to_signed(0, 8), to_signed(180, 8), to_signed(180, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(201, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(173, 8), to_signed(173, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(118, 8), to_signed(118, 8), to_signed(40, 8), to_signed(0, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(45, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(173, 8), to_signed(173, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(85, 8), to_signed(118, 8), to_signed(85, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(201, 8), 
to_signed(40, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(173, 8), to_signed(173, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(45, 8), 
to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(201, 8), 
to_signed(40, 8), to_signed(28, 8), to_signed(0, 8), to_signed(85, 8), to_signed(85, 8), to_signed(45, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(173, 8), to_signed(173, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(45, 8), to_signed(173, 8), to_signed(173, 8), 
to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(201, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(85, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(45, 8), to_signed(173, 8), to_signed(173, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(85, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(0, 8), to_signed(8, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(44, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(0, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(48, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(44, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(44, 8), to_signed(8, 8), to_signed(44, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(72, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(104, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(218, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(73, 8), to_signed(218, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(73, 8), to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(73, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(218, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(218, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(73, 8), to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(72, 8), to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(77, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(140, 8), to_signed(72, 8), to_signed(72, 8), to_signed(72, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(218, 8), to_signed(73, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(77, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), 
to_signed(218, 8), to_signed(145, 8), to_signed(77, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(72, 8), to_signed(104, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(72, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(218, 8), to_signed(73, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(218, 8), to_signed(182, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(73, 8), to_signed(73, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(77, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(0, 8), to_signed(145, 8), to_signed(218, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(77, 8), to_signed(145, 8), to_signed(0, 8), to_signed(0, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(77, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(140, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(72, 8), to_signed(72, 8), to_signed(72, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(182, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(73, 8), to_signed(145, 8), to_signed(0, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(140, 8), to_signed(72, 8), to_signed(104, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(73, 8), to_signed(145, 8), to_signed(145, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(145, 8), to_signed(145, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(73, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(48, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(77, 8), to_signed(145, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(73, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(77, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(104, 8), to_signed(72, 8), to_signed(0, 8), 
to_signed(8, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(77, 8), to_signed(145, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(77, 8), 
to_signed(73, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(77, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(77, 8), to_signed(145, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(77, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(73, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(145, 8), to_signed(0, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(73, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(145, 8), to_signed(77, 8), to_signed(73, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(145, 8), to_signed(73, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(145, 8), to_signed(77, 8), to_signed(0, 8), to_signed(0, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(77, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(77, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(48, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(77, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(218, 8), to_signed(77, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(73, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(218, 8), to_signed(77, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(73, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(218, 8), to_signed(145, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(8, 8), to_signed(48, 8), to_signed(218, 8), to_signed(145, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(77, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(145, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(48, 8), to_signed(8, 8), to_signed(48, 8), to_signed(0, 8), to_signed(218, 8), to_signed(145, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(8, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(77, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(218, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(77, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(73, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(73, 8), to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(73, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(77, 8), to_signed(145, 8), to_signed(77, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(73, 8), 
to_signed(145, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(77, 8), to_signed(73, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(0, 8), to_signed(76, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(73, 8), to_signed(77, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(77, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(76, 8), to_signed(76, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(28, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(8, 8), to_signed(48, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(44, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), 
to_signed(48, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(48, 8), 
to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(44, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(145, 8), to_signed(218, 8), to_signed(182, 8), to_signed(77, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(8, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(145, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(72, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(145, 8), to_signed(218, 8), to_signed(145, 8), to_signed(182, 8), to_signed(77, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(72, 8), to_signed(0, 8), to_signed(72, 8), to_signed(72, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(145, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(72, 8), to_signed(72, 8), to_signed(72, 8), 
to_signed(72, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(48, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(44, 8), to_signed(48, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(8, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(145, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(182, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(72, 8), 
to_signed(72, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(44, 8), to_signed(48, 8), to_signed(44, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(77, 8), to_signed(182, 8), to_signed(182, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(44, 8), 
to_signed(0, 8), to_signed(72, 8), to_signed(104, 8), to_signed(0, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(77, 8), to_signed(77, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), to_signed(182, 8), to_signed(182, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(0, 8), to_signed(77, 8), to_signed(182, 8), to_signed(182, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(72, 8), 
to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(77, 8), to_signed(182, 8), to_signed(77, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(8, 8), 
to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(8, 8), to_signed(72, 8), to_signed(72, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(72, 8), to_signed(0, 8), to_signed(44, 8), to_signed(44, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(44, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(77, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), 
to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(44, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), 
to_signed(72, 8), to_signed(72, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(77, 8), to_signed(28, 8), to_signed(28, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(182, 8), to_signed(182, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(77, 8), 
to_signed(77, 8), to_signed(77, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(0, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(40, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(0, 8), to_signed(72, 8), to_signed(72, 8), to_signed(72, 8), to_signed(72, 8), to_signed(28, 8), to_signed(72, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(0, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(40, 8), 
to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(72, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(104, 8), to_signed(0, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), 
to_signed(8, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(72, 8), to_signed(72, 8), to_signed(140, 8), to_signed(72, 8), to_signed(72, 8), to_signed(72, 8), to_signed(72, 8), 
to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(8, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(8, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(44, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(72, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(140, 8), to_signed(72, 8), to_signed(104, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(104, 8), to_signed(72, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(48, 8), to_signed(44, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), to_signed(72, 8), to_signed(140, 8), to_signed(72, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(8, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(72, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(145, 8), to_signed(72, 8), to_signed(72, 8), to_signed(8, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(8, 8), to_signed(140, 8), to_signed(140, 8), to_signed(72, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(40, 8), to_signed(145, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(145, 8), to_signed(145, 8), to_signed(145, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(72, 8), to_signed(140, 8), to_signed(104, 8), to_signed(72, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(40, 8), to_signed(145, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), to_signed(145, 8), 
to_signed(145, 8), to_signed(40, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(44, 8), 
to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(44, 8), to_signed(72, 8), to_signed(140, 8), to_signed(104, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(145, 8), to_signed(145, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(0, 8), to_signed(72, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(72, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(40, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(48, 8), to_signed(48, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(72, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(40, 8), to_signed(76, 8), to_signed(76, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(40, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), 
to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(40, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(40, 8), to_signed(40, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(76, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(76, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(104, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(182, 8), to_signed(0, 8), to_signed(40, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(40, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(218, 8), to_signed(77, 8), to_signed(0, 8), to_signed(0, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(76, 8), to_signed(40, 8), to_signed(76, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(76, 8), to_signed(76, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(104, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(104, 8), to_signed(218, 8), to_signed(182, 8), to_signed(0, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(77, 8), to_signed(73, 8), to_signed(0, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(76, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(76, 8), to_signed(76, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(40, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(0, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(40, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(0, 8), to_signed(76, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(40, 8), to_signed(76, 8), to_signed(104, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(40, 8), to_signed(48, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(76, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(76, 8), to_signed(76, 8), to_signed(0, 8), to_signed(76, 8), to_signed(76, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(40, 8), to_signed(76, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(40, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(76, 8), to_signed(73, 8), to_signed(73, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(76, 8), to_signed(140, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(182, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(40, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(73, 8), to_signed(73, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(40, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(40, 8), to_signed(72, 8), to_signed(72, 8), to_signed(76, 8), to_signed(76, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(140, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(0, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(73, 8), to_signed(104, 8), to_signed(0, 8), to_signed(48, 8), to_signed(76, 8), to_signed(40, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(73, 8), to_signed(73, 8), to_signed(48, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(40, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(72, 8), to_signed(72, 8), to_signed(104, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(140, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(0, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), 
to_signed(76, 8), to_signed(73, 8), to_signed(218, 8), to_signed(218, 8), to_signed(0, 8), to_signed(76, 8), to_signed(76, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(73, 8), to_signed(48, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(40, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(72, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(48, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(76, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(73, 8), to_signed(182, 8), to_signed(73, 8), to_signed(72, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(48, 8), to_signed(48, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(40, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(77, 8), to_signed(73, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(0, 8), to_signed(0, 8), to_signed(140, 8), to_signed(72, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(48, 8), to_signed(72, 8), to_signed(72, 8), to_signed(72, 8), 
to_signed(72, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(40, 8), to_signed(76, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(0, 8), to_signed(73, 8), to_signed(77, 8), to_signed(77, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(72, 8), to_signed(40, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), 
to_signed(40, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(76, 8), to_signed(48, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(104, 8), to_signed(72, 8), to_signed(76, 8), to_signed(72, 8), to_signed(40, 8), to_signed(72, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(72, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(73, 8), to_signed(0, 8), 
to_signed(72, 8), to_signed(72, 8), to_signed(72, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(40, 8), to_signed(40, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(0, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(72, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), 
to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(76, 8), to_signed(0, 8), to_signed(72, 8), to_signed(72, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(72, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(40, 8), 
to_signed(40, 8), to_signed(40, 8), to_signed(0, 8), to_signed(0, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(72, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(72, 8), to_signed(140, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(72, 8), 
to_signed(72, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(72, 8), to_signed(140, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(72, 8), 
to_signed(72, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(72, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(72, 8), to_signed(140, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(72, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(72, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(72, 8), to_signed(182, 8), 
to_signed(77, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(72, 8), to_signed(140, 8), to_signed(72, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(72, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(104, 8), to_signed(72, 8), to_signed(104, 8), to_signed(72, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(72, 8), to_signed(72, 8), to_signed(72, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(73, 8), to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(72, 8), to_signed(182, 8), to_signed(104, 8), to_signed(72, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(72, 8), to_signed(182, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(73, 8), to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(73, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(72, 8), to_signed(182, 8), to_signed(72, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(73, 8), to_signed(182, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(104, 8), to_signed(72, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(72, 8), to_signed(104, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(140, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(104, 8), to_signed(72, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(72, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), 
to_signed(77, 8), to_signed(218, 8), to_signed(77, 8), to_signed(104, 8), to_signed(104, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(77, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(104, 8), to_signed(140, 8), to_signed(140, 8), to_signed(104, 8), to_signed(77, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(77, 8), to_signed(182, 8), to_signed(72, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), to_signed(104, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(218, 8), to_signed(104, 8), to_signed(104, 8), to_signed(77, 8), to_signed(218, 8), 
to_signed(218, 8), to_signed(218, 8), to_signed(218, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(73, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(132, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(168, 8), to_signed(132, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(204, 8), to_signed(132, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(141, 8), to_signed(141, 8), to_signed(141, 8), to_signed(109, 8), to_signed(109, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(132, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(141, 8), to_signed(141, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(204, 8), to_signed(204, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(141, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(204, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(109, 8), to_signed(141, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(36, 8), to_signed(132, 8), to_signed(204, 8), 
to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(141, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(204, 8), to_signed(168, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(141, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(109, 8), to_signed(141, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), 
to_signed(141, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(141, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(141, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), 
to_signed(141, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(141, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(141, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(177, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(141, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(177, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(177, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(109, 8), to_signed(177, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), 
to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(177, 8), to_signed(109, 8), to_signed(109, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(177, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(109, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(177, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(177, 8), to_signed(0, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(109, 8), to_signed(109, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(36, 8), to_signed(0, 8), to_signed(168, 8), to_signed(0, 8), to_signed(177, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(178, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(177, 8), to_signed(36, 8), 
to_signed(0, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(177, 8), 
to_signed(0, 8), to_signed(177, 8), to_signed(0, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(178, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(109, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(177, 8), to_signed(36, 8), to_signed(0, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(0, 8), to_signed(217, 8), to_signed(213, 8), to_signed(0, 8), 
to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(178, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(109, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(177, 8), to_signed(177, 8), to_signed(36, 8), to_signed(0, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(217, 8), to_signed(109, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(109, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(177, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(36, 8), to_signed(0, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(217, 8), to_signed(0, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(109, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(177, 8), to_signed(36, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(177, 8), to_signed(177, 8), 
to_signed(213, 8), to_signed(177, 8), to_signed(177, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(109, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(177, 8), to_signed(109, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(177, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(132, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(177, 8), to_signed(177, 8), to_signed(0, 8), 
to_signed(177, 8), to_signed(213, 8), to_signed(177, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(178, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(109, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(177, 8), to_signed(177, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(132, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(132, 8), to_signed(178, 8), to_signed(109, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(213, 8), to_signed(177, 8), to_signed(109, 8), to_signed(177, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(109, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(177, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), 
to_signed(178, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(177, 8), to_signed(109, 8), to_signed(36, 8), to_signed(177, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(109, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(109, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), 
to_signed(178, 8), to_signed(109, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(178, 8), to_signed(178, 8), to_signed(0, 8), 
to_signed(213, 8), to_signed(36, 8), to_signed(168, 8), to_signed(36, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(109, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(0, 8), to_signed(109, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), 
to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), to_signed(0, 8), to_signed(178, 8), to_signed(178, 8), to_signed(0, 8), to_signed(168, 8), 
to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(109, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(0, 8), to_signed(204, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(109, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(213, 8), to_signed(109, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(0, 8), to_signed(109, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(0, 8), to_signed(109, 8), 
to_signed(213, 8), to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), to_signed(0, 8), to_signed(204, 8), to_signed(168, 8), 
to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(36, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(109, 8), to_signed(178, 8), to_signed(213, 8), to_signed(36, 8), to_signed(0, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(168, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(36, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), to_signed(213, 8), 
to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(36, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(168, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(36, 8), 
to_signed(109, 8), to_signed(36, 8), to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), 
to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(109, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), 
to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), 
to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), 
to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), to_signed(109, 8), 
to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(168, 8), to_signed(168, 8), to_signed(132, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(109, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(109, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(168, 8), to_signed(132, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(132, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(36, 8), to_signed(0, 8), to_signed(36, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(132, 8), to_signed(168, 8), to_signed(132, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(132, 8), to_signed(168, 8), to_signed(132, 8), to_signed(132, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(168, 8), to_signed(168, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(132, 8), to_signed(132, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(132, 8), to_signed(168, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(132, 8), to_signed(168, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(132, 8), to_signed(168, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(132, 8), to_signed(168, 8), to_signed(168, 8), to_signed(132, 8), to_signed(168, 8), to_signed(132, 8), to_signed(168, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(132, 8), to_signed(168, 8), to_signed(132, 8), to_signed(168, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(109, 8), to_signed(204, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(213, 8), to_signed(177, 8), to_signed(213, 8), to_signed(177, 8), to_signed(204, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(168, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), 
to_signed(177, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(204, 8), to_signed(132, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(204, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(213, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(177, 8), to_signed(204, 8), to_signed(36, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(204, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(204, 8), to_signed(204, 8), to_signed(36, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(204, 8), to_signed(36, 8), to_signed(28, 8), to_signed(177, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(177, 8), to_signed(204, 8), to_signed(132, 8), to_signed(213, 8), to_signed(213, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(36, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(204, 8), to_signed(36, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(213, 8), to_signed(204, 8), to_signed(204, 8), to_signed(36, 8), to_signed(177, 8), to_signed(36, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), 
to_signed(217, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(141, 8), to_signed(204, 8), to_signed(132, 8), to_signed(36, 8), to_signed(0, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(204, 8), to_signed(168, 8), to_signed(36, 8), to_signed(0, 8), to_signed(213, 8), to_signed(132, 8), to_signed(168, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(168, 8), to_signed(204, 8), to_signed(36, 8), 
to_signed(109, 8), to_signed(204, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(213, 8), to_signed(132, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(177, 8), to_signed(213, 8), to_signed(141, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(36, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(204, 8), to_signed(132, 8), 
to_signed(204, 8), to_signed(168, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(141, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(168, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(168, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(132, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(141, 8), to_signed(141, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(213, 8), 
to_signed(204, 8), to_signed(132, 8), to_signed(132, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(36, 8), to_signed(36, 8), to_signed(177, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(217, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(132, 8), to_signed(132, 8), to_signed(36, 8), to_signed(36, 8), to_signed(168, 8), to_signed(36, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(36, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(168, 8), to_signed(0, 8), to_signed(0, 8), to_signed(132, 8), to_signed(132, 8), to_signed(36, 8), to_signed(177, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(177, 8), to_signed(213, 8), to_signed(132, 8), to_signed(168, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(168, 8), to_signed(36, 8), to_signed(178, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(141, 8), to_signed(141, 8), to_signed(36, 8), to_signed(109, 8), to_signed(109, 8), to_signed(177, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(213, 8), to_signed(132, 8), to_signed(132, 8), to_signed(168, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), to_signed(36, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(141, 8), to_signed(141, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(177, 8), to_signed(213, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(132, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), to_signed(36, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(141, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(109, 8), to_signed(213, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(132, 8), to_signed(132, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), 
to_signed(141, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(0, 8), to_signed(0, 8), to_signed(177, 8), 
to_signed(0, 8), to_signed(36, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), 
to_signed(36, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(109, 8), to_signed(141, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(36, 8), to_signed(36, 8), to_signed(217, 8), to_signed(213, 8), to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(178, 8), to_signed(177, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(109, 8), to_signed(0, 8), to_signed(168, 8), to_signed(204, 8), to_signed(204, 8), to_signed(109, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(36, 8), to_signed(109, 8), to_signed(109, 8), to_signed(141, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(213, 8), to_signed(36, 8), 
to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(177, 8), to_signed(177, 8), 
to_signed(177, 8), to_signed(177, 8), to_signed(0, 8), to_signed(0, 8), to_signed(204, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(141, 8), to_signed(213, 8), to_signed(36, 8), to_signed(177, 8), to_signed(177, 8), to_signed(109, 8), to_signed(109, 8), to_signed(141, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(217, 8), to_signed(213, 8), to_signed(109, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(36, 8), to_signed(177, 8), to_signed(213, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), 
to_signed(109, 8), to_signed(0, 8), to_signed(109, 8), to_signed(109, 8), to_signed(0, 8), to_signed(109, 8), to_signed(178, 8), to_signed(141, 8), 
to_signed(213, 8), to_signed(141, 8), to_signed(141, 8), to_signed(36, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), 
to_signed(109, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(109, 8), to_signed(132, 8), to_signed(204, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(132, 8), to_signed(36, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(109, 8), to_signed(109, 8), to_signed(36, 8), to_signed(141, 8), 
to_signed(178, 8), to_signed(178, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(177, 8), to_signed(177, 8), to_signed(177, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(177, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(178, 8), 
to_signed(178, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(109, 8), to_signed(217, 8), to_signed(213, 8), to_signed(178, 8), to_signed(109, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(132, 8), to_signed(36, 8), to_signed(177, 8), to_signed(109, 8), to_signed(177, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), to_signed(213, 8), to_signed(178, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(213, 8), to_signed(178, 8), 
to_signed(0, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), 
to_signed(178, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(109, 8), to_signed(217, 8), to_signed(109, 8), to_signed(178, 8), to_signed(109, 8), to_signed(132, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(36, 8), to_signed(178, 8), to_signed(213, 8), to_signed(178, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(109, 8), to_signed(109, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(217, 8), to_signed(178, 8), to_signed(178, 8), 
to_signed(141, 8), to_signed(36, 8), to_signed(36, 8), to_signed(109, 8), to_signed(178, 8), to_signed(109, 8), to_signed(178, 8), to_signed(0, 8), 
to_signed(109, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(28, 8), to_signed(109, 8), to_signed(0, 8), to_signed(132, 8), to_signed(132, 8), 
to_signed(209, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(141, 8), to_signed(109, 8), to_signed(141, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(178, 8), to_signed(178, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(217, 8), to_signed(36, 8), to_signed(141, 8), 
to_signed(141, 8), to_signed(109, 8), to_signed(141, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(168, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(168, 8), to_signed(132, 8), to_signed(0, 8), to_signed(132, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(109, 8), to_signed(217, 8), to_signed(109, 8), to_signed(0, 8), to_signed(141, 8), to_signed(36, 8), 
to_signed(141, 8), to_signed(109, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(141, 8), to_signed(109, 8), to_signed(178, 8), to_signed(178, 8), to_signed(178, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(204, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(132, 8), to_signed(132, 8), to_signed(168, 8), to_signed(132, 8), to_signed(168, 8), to_signed(36, 8), to_signed(132, 8), 
to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(217, 8), to_signed(0, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(36, 8), to_signed(217, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(141, 8), to_signed(141, 8), to_signed(141, 8), 
to_signed(141, 8), to_signed(141, 8), to_signed(109, 8), to_signed(141, 8), to_signed(178, 8), to_signed(178, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(109, 8), to_signed(0, 8), to_signed(217, 8), to_signed(0, 8), to_signed(109, 8), to_signed(109, 8), to_signed(36, 8), 
to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(141, 8), to_signed(141, 8), to_signed(141, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(141, 8), to_signed(141, 8), to_signed(141, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(168, 8), to_signed(36, 8), to_signed(132, 8), to_signed(132, 8), to_signed(132, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), to_signed(0, 8), to_signed(109, 8), to_signed(36, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(178, 8), to_signed(178, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(109, 8), to_signed(141, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(168, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(141, 8), to_signed(109, 8), to_signed(109, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(109, 8), 
to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(178, 8), to_signed(178, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(168, 8), to_signed(204, 8), to_signed(204, 8), to_signed(132, 8), to_signed(168, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(217, 8), to_signed(217, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(204, 8), to_signed(204, 8), to_signed(132, 8), to_signed(36, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(168, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(109, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(36, 8), to_signed(132, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(36, 8), 
to_signed(168, 8), to_signed(36, 8), to_signed(168, 8), to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(168, 8), to_signed(132, 8), to_signed(168, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(168, 8), to_signed(0, 8), to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(28, 8), to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(168, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(132, 8), to_signed(204, 8), to_signed(204, 8), to_signed(209, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(168, 8), to_signed(204, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(132, 8), to_signed(168, 8), to_signed(204, 8), to_signed(213, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(168, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(209, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(168, 8), to_signed(209, 8), to_signed(213, 8), to_signed(209, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(168, 8), 
to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(204, 8), to_signed(213, 8), to_signed(204, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(168, 8), to_signed(209, 8), to_signed(213, 8), to_signed(209, 8), to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(204, 8), to_signed(204, 8), to_signed(168, 8), to_signed(213, 8), to_signed(209, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(168, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(209, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(209, 8), to_signed(213, 8), to_signed(209, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(209, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), to_signed(168, 8), to_signed(168, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(168, 8), to_signed(209, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), to_signed(168, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(132, 8), 
to_signed(209, 8), to_signed(168, 8), to_signed(168, 8), to_signed(209, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), to_signed(168, 8), 
to_signed(168, 8), to_signed(209, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), 
to_signed(213, 8), to_signed(168, 8), to_signed(168, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), 
to_signed(168, 8), to_signed(209, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), 
to_signed(213, 8), to_signed(209, 8), to_signed(168, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), 
to_signed(168, 8), to_signed(209, 8), to_signed(209, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), 
to_signed(209, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), 
to_signed(213, 8), to_signed(209, 8), to_signed(209, 8), to_signed(109, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(168, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(109, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(209, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), 
to_signed(213, 8), to_signed(209, 8), to_signed(209, 8), to_signed(109, 8), to_signed(209, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(109, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(109, 8), to_signed(209, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), to_signed(209, 8), 
to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), 
to_signed(109, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), 
to_signed(36, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(209, 8), to_signed(209, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), to_signed(0, 8), to_signed(213, 8), to_signed(213, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(213, 8), 
to_signed(36, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), to_signed(109, 8), to_signed(109, 8), to_signed(209, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(109, 8), to_signed(109, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), 
to_signed(213, 8), to_signed(213, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(109, 8), to_signed(213, 8), to_signed(36, 8), to_signed(36, 8), to_signed(213, 8), to_signed(213, 8), to_signed(213, 8), to_signed(109, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(109, 8), to_signed(209, 8), to_signed(209, 8), to_signed(209, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(213, 8), to_signed(213, 8), to_signed(36, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(68, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(136, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(136, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(216, 8), to_signed(212, 8), 
to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(216, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(136, 8), to_signed(212, 8), to_signed(68, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), 
to_signed(68, 8), to_signed(36, 8), to_signed(36, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(68, 8), to_signed(136, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(36, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(136, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(68, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(208, 8), 
to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(68, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(136, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(136, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(68, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), 
to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(208, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(208, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(208, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(200, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(200, 8), to_signed(160, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(160, 8), to_signed(160, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(68, 8), to_signed(208, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(160, 8), to_signed(160, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(36, 8), to_signed(208, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(160, 8), to_signed(160, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(200, 8), to_signed(160, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(136, 8), to_signed(208, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(208, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(136, 8), to_signed(208, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(208, 8), to_signed(36, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(208, 8), to_signed(36, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(208, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(36, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(36, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), 
to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(208, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(208, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(68, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(36, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(36, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(136, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(212, 8), to_signed(208, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(208, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(208, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(36, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(208, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), 
to_signed(68, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(36, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(136, 8), to_signed(212, 8), to_signed(136, 8), to_signed(212, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), 
to_signed(68, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(68, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(36, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(68, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(36, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(68, 8), to_signed(36, 8), to_signed(68, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(136, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(208, 8), to_signed(208, 8), to_signed(36, 8), to_signed(36, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(208, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(36, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(136, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(36, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(36, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(208, 8), to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(136, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(212, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(136, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(136, 8), to_signed(208, 8), to_signed(249, 8), to_signed(249, 8), 
to_signed(249, 8), to_signed(216, 8), to_signed(216, 8), to_signed(208, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(208, 8), to_signed(249, 8), to_signed(249, 8), to_signed(249, 8), to_signed(249, 8), 
to_signed(249, 8), to_signed(249, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(68, 8), to_signed(208, 8), to_signed(216, 8), to_signed(249, 8), to_signed(249, 8), to_signed(249, 8), to_signed(249, 8), to_signed(249, 8), 
to_signed(249, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(208, 8), 
to_signed(136, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(208, 8), to_signed(0, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(73, 8), to_signed(255, 8), to_signed(0, 8), to_signed(36, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(0, 8), to_signed(255, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(36, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), to_signed(68, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(208, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), 
to_signed(36, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(200, 8), to_signed(200, 8), to_signed(216, 8), 
to_signed(208, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(68, 8), to_signed(136, 8), to_signed(208, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(160, 8), 
to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(200, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(208, 8), to_signed(68, 8), to_signed(136, 8), to_signed(160, 8), to_signed(160, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(208, 8), to_signed(216, 8), to_signed(212, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), 
to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(160, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), 
to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), to_signed(160, 8), 
to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(160, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(200, 8), to_signed(200, 8), 
to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(160, 8), to_signed(160, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(200, 8), to_signed(200, 8), 
to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(136, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(208, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(208, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(0, 8), to_signed(68, 8), to_signed(208, 8), to_signed(208, 8), to_signed(208, 8), 
to_signed(212, 8), to_signed(208, 8), to_signed(68, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(208, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(0, 8), to_signed(208, 8), to_signed(208, 8), to_signed(208, 8), to_signed(208, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(208, 8), to_signed(208, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(0, 8), to_signed(208, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(208, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(0, 8), to_signed(216, 8), to_signed(208, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(136, 8), to_signed(136, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(136, 8), to_signed(136, 8), 
to_signed(136, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(68, 8), to_signed(136, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(216, 8), to_signed(212, 8), 
to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), to_signed(216, 8), 
to_signed(216, 8), to_signed(216, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(216, 8), to_signed(212, 8), to_signed(216, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(136, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(208, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(68, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(208, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(208, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(136, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(68, 8), to_signed(136, 8), to_signed(136, 8), to_signed(208, 8), 
to_signed(208, 8), to_signed(136, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(216, 8), to_signed(136, 8), 
to_signed(216, 8), to_signed(208, 8), to_signed(68, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(136, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(216, 8), to_signed(136, 8), to_signed(216, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(138, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(138, 8), to_signed(174, 8), to_signed(101, 8), to_signed(101, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(174, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(68, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(138, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(101, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(101, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(28, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(28, 8), 
to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(68, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(68, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(68, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(68, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(174, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(174, 8), to_signed(174, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(0, 8), to_signed(138, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(68, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(0, 8), to_signed(174, 8), to_signed(174, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(68, 8), to_signed(0, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(0, 8), to_signed(68, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(0, 8), to_signed(164, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(174, 8), to_signed(0, 8), to_signed(164, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(241, 8), to_signed(68, 8), to_signed(138, 8), to_signed(174, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(241, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(241, 8), to_signed(164, 8), to_signed(0, 8), to_signed(138, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(200, 8), to_signed(200, 8), to_signed(0, 8), to_signed(101, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(68, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(68, 8), to_signed(28, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(164, 8), to_signed(200, 8), to_signed(164, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(164, 8), to_signed(68, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(214, 8), to_signed(68, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), to_signed(68, 8), to_signed(0, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(214, 8), 
to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(68, 8), to_signed(138, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(68, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(214, 8), to_signed(73, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(251, 8), to_signed(251, 8), to_signed(73, 8), to_signed(214, 8), to_signed(214, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(251, 8), to_signed(251, 8), to_signed(73, 8), to_signed(251, 8), to_signed(214, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(251, 8), to_signed(214, 8), to_signed(251, 8), to_signed(73, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(68, 8), to_signed(251, 8), to_signed(214, 8), to_signed(73, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(68, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(251, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(0, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(68, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(101, 8), to_signed(138, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(68, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(174, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(101, 8), to_signed(138, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(138, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(101, 8), to_signed(174, 8), to_signed(101, 8), to_signed(28, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(28, 8), to_signed(101, 8), to_signed(138, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(101, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(101, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(174, 8), to_signed(138, 8), 
to_signed(68, 8), to_signed(101, 8), to_signed(174, 8), to_signed(138, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), 
to_signed(101, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(138, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(138, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(68, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(138, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(174, 8), to_signed(138, 8), to_signed(174, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(101, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(68, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(68, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(68, 8), to_signed(138, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(200, 8), to_signed(200, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(138, 8), to_signed(68, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(174, 8), to_signed(138, 8), to_signed(68, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(0, 8), to_signed(0, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(200, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(174, 8), to_signed(174, 8), 
to_signed(138, 8), to_signed(0, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(68, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(200, 8), to_signed(200, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(174, 8), to_signed(138, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(0, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(200, 8), to_signed(0, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(164, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(0, 8), to_signed(200, 8), 
to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(0, 8), 
to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(101, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(164, 8), to_signed(200, 8), to_signed(200, 8), to_signed(200, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), 
to_signed(214, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(200, 8), to_signed(200, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(68, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(68, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(68, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(251, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(68, 8), to_signed(68, 8), to_signed(73, 8), to_signed(214, 8), to_signed(251, 8), to_signed(251, 8), to_signed(214, 8), 
to_signed(68, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(0, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(251, 8), to_signed(73, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(73, 8), to_signed(214, 8), to_signed(214, 8), to_signed(73, 8), to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(68, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(214, 8), to_signed(73, 8), to_signed(214, 8), to_signed(214, 8), 
to_signed(214, 8), to_signed(73, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(214, 8), to_signed(73, 8), to_signed(251, 8), 
to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(178, 8), to_signed(178, 8), to_signed(251, 8), to_signed(214, 8), to_signed(68, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(73, 8), to_signed(251, 8), to_signed(251, 8), 
to_signed(251, 8), to_signed(73, 8), to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(73, 8), to_signed(251, 8), 
to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(73, 8), to_signed(251, 8), to_signed(68, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(251, 8), to_signed(251, 8), 
to_signed(251, 8), to_signed(178, 8), to_signed(178, 8), to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(178, 8), to_signed(178, 8), 
to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(73, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(251, 8), 
to_signed(251, 8), to_signed(251, 8), to_signed(73, 8), to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(73, 8), 
to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(68, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(251, 8), to_signed(73, 8), to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(251, 8), to_signed(73, 8), 
to_signed(251, 8), to_signed(68, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), to_signed(68, 8), 
to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(138, 8), to_signed(68, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(68, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(101, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(68, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), 
to_signed(68, 8), to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(68, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(68, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(174, 8), to_signed(174, 8), to_signed(174, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(68, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(138, 8), to_signed(174, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(68, 8), to_signed(0, 8), to_signed(68, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(138, 8), to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(68, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(68, 8), to_signed(68, 8), to_signed(138, 8), 
to_signed(138, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(101, 8), 
to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(0, 8), to_signed(101, 8), to_signed(101, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(46, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), to_signed(82, 8), to_signed(46, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(46, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(82, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), to_signed(82, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(77, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(82, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(255, 8), to_signed(0, 8), to_signed(77, 8), to_signed(255, 8), 
to_signed(82, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(255, 8), to_signed(0, 8), to_signed(0, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(77, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), 
to_signed(255, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(77, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(0, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(77, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(77, 8), to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(0, 8), to_signed(0, 8), to_signed(77, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(77, 8), to_signed(212, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), to_signed(77, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(140, 8), to_signed(72, 8), to_signed(72, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(77, 8), to_signed(140, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(77, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(182, 8), to_signed(182, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(82, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(46, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(0, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), to_signed(9, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(9, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), 
to_signed(46, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(46, 8), to_signed(46, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(82, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(150, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(182, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(182, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(150, 8), to_signed(46, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(46, 8), to_signed(82, 8), to_signed(150, 8), to_signed(9, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(255, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(82, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(182, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(255, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(82, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(255, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(150, 8), to_signed(82, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(182, 8), to_signed(77, 8), 
to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(182, 8), to_signed(82, 8), to_signed(150, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(150, 8), to_signed(82, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(0, 8), to_signed(255, 8), 
to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(182, 8), to_signed(182, 8), to_signed(140, 8), to_signed(250, 8), 
to_signed(250, 8), to_signed(82, 8), to_signed(82, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(0, 8), to_signed(255, 8), 
to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(140, 8), to_signed(250, 8), to_signed(250, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(140, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(140, 8), to_signed(250, 8), to_signed(212, 8), 
to_signed(212, 8), to_signed(212, 8), to_signed(72, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(77, 8), to_signed(0, 8), 
to_signed(77, 8), to_signed(255, 8), to_signed(255, 8), to_signed(182, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(77, 8), to_signed(72, 8), to_signed(212, 8), 
to_signed(140, 8), to_signed(72, 8), to_signed(140, 8), to_signed(182, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(72, 8), 
to_signed(72, 8), to_signed(140, 8), to_signed(72, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(182, 8), to_signed(182, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), to_signed(182, 8), 
to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(46, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(46, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(46, 8), to_signed(9, 8), to_signed(0, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(0, 8), to_signed(46, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(150, 8), to_signed(9, 8), to_signed(46, 8), 
to_signed(46, 8), to_signed(9, 8), to_signed(0, 8), to_signed(150, 8), to_signed(150, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(9, 8), to_signed(46, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), 
to_signed(150, 8), to_signed(82, 8), to_signed(9, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(82, 8), to_signed(9, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(82, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(9, 8), to_signed(255, 8), to_signed(182, 8), to_signed(150, 8), to_signed(150, 8), to_signed(182, 8), to_signed(255, 8), 
to_signed(182, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(9, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(150, 8), 
to_signed(150, 8), to_signed(9, 8), to_signed(255, 8), to_signed(255, 8), to_signed(150, 8), to_signed(150, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(9, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(82, 8), to_signed(255, 8), to_signed(150, 8), to_signed(150, 8), to_signed(182, 8), to_signed(255, 8), 
to_signed(182, 8), to_signed(150, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), to_signed(82, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(150, 8), to_signed(150, 8), to_signed(150, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(150, 8), to_signed(150, 8), to_signed(9, 8), to_signed(82, 8), to_signed(9, 8), 
to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), 
to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(140, 8), to_signed(72, 8), to_signed(72, 8), to_signed(140, 8), to_signed(140, 8), to_signed(140, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(9, 8), to_signed(82, 8), to_signed(82, 8), to_signed(82, 8), to_signed(9, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(72, 8), to_signed(212, 8), to_signed(140, 8), to_signed(212, 8), to_signed(140, 8), to_signed(72, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(9, 8), to_signed(9, 8), to_signed(140, 8), to_signed(140, 8), to_signed(72, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(72, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(140, 8), to_signed(212, 8), to_signed(212, 8), to_signed(140, 8), to_signed(0, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(140, 8), to_signed(250, 8), to_signed(140, 8), to_signed(250, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8));