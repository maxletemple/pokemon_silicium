type rom_type is array (0 TO 2394) of signed (7 DOWNTO 0);
signal rom : rom_type := (to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(146, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(146, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(0, 8), to_signed(146, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(146, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), 
to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(255, 8), to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), to_signed(146, 8), 
to_signed(146, 8), to_signed(146, 8), to_signed(0, 8), to_signed(0, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), to_signed(28, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(28, 8), to_signed(28, 8), to_signed(0, 8));