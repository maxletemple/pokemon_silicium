LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY rom_arenas IS
    PORT (
        CLOCK          : IN  STD_LOGIC;
        ADDR_R         : IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
        DATA_OUT       : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END rom_arenas;

ARCHITECTURE Behavioral OF rom_arenas IS
    type rom_type is array (0 TO 28160) of signed (7 DOWNTO 0);
signal rom : rom_type := (to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), 
to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(37, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(4, 8), to_signed(1, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(41, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(41, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), to_signed(41, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), 
to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(41, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(37, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(5, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), 
to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(4, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(0, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(0, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(37, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(37, 8), to_signed(37, 8), to_signed(5, 8), to_signed(37, 8), to_signed(37, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(0, 8), to_signed(1, 8), to_signed(0, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(0, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(1, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(36, 8), to_signed(73, 8), to_signed(69, 8), to_signed(73, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(0, 8), to_signed(0, 8), to_signed(0, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(36, 8), 
to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(69, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(69, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(69, 8), to_signed(69, 8), 
to_signed(73, 8), to_signed(73, 8), to_signed(73, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), 
to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(36, 8), to_signed(0, 8), 
to_signed(0, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), 
to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(5, 8), to_signed(5, 8), to_signed(5, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), to_signed(1, 8), 
to_signed(0, 8));
    -- QUELQUES PETITES MODIFICATIONS FAITES POUR AIDER VIVADO A FAIRE LES BONS
    -- CHOIX D'IMPLEMENTATION...

    ATTRIBUTE RAM_STYLE : string;
    ATTRIBUTE RAM_STYLE of rom: signal is "BLOCK";

BEGIN

    PROCESS (CLOCK)
    BEGIN
        IF (CLOCK'event AND CLOCK = '1') THEN
            if (unsigned(addr_r) <= to_unsigned(28160, 16)) then
                DATA_OUT <= STD_LOGIC_VECTOR( rom(to_integer(UNSIGNED(ADDR_R))) );
            end if;
        END IF;
    END PROCESS;

END Behavioral;