LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY rom_letters IS
PORT (
      CLOCK          : IN  STD_LOGIC;
      ADDR_R         : IN  STD_LOGIC_VECTOR(6 DOWNTO 0);
      DATA_OUT       : OUT STD_LOGIC_VECTOR(39 DOWNTO 0)
      );
END rom_letters;

ARCHITECTURE Behavioral OF rom_letters IS
type rom_type is array (0 TO 78) of std_logic_vector (39 DOWNTO 0);
signal rom : rom_type := ("0110010010100101111010010100101001000000", "1110010010100101110010010100101110000000", "0110010010100001000010000100100110000000", "1110010010100101001010010100101110000000", "1111010000100001110010000100001111000000", "1111010000100001110010000100001000000000", "0110010010100001011010010100100110000000", "1001010010100101111010010100101001000000", "1110001000010000100001000010001110000000", "0001000010000100001010010100100110000000", "1001010010101001100010100100101001000000", "1000010000100001000010000100001111000000", "1001011110100101001010010100101001000000", "1001011010110101011010110100101001000000", "0110010010100101001010010100100110000000", "1110010010100101110010000100001000000000", "0110010010100101001010010101100110000010", "1110010010100101110010010100101001000000", "0110010010100000110000010100100110000000", "0111000100001000010000100001000010000000", "1001010010100101001010010100100110000000", "1001010010100101001010010101000100000000", "1001010010100101001010010111101001000000", "1001010010100100110010010100101001000000", "1010010100101001010001000010000100000000", "1111000010001000010001000010001111000000", "0000000000011101001010010101100101000000", "1000010000111001001010010100101110000000", "0000000000011001001010000100100110000000", "0001000010011101001010010100100111000000", "0000000000011001001011110100000111000000", "0011001000111000100001000010000100000000", "0000001110100101001001110000100110000000", "1000010000111001001010010100101001000000", "0010000000001000010000100001000010000000", "0010000000001000010000100001001100000000", "1000010000100101010011000101001001000000", "0010000100001000010000100001000010000000", "0000000000110111010110101101011010100000", "0000000000111001001010010100101001000000", "0000000000011001001010010100100110000000", "0000000000111001001010010111001000010000", "0000000000011101001010010011100001000010", "0000000000101101100010000100001000000000", "0000000000011101000001100000101110000000", "0000001000111100100001000010000011000000", "0000000000100101001010010101100101000000", "0000000000100101001010010101000100000000", "0000000000100101001010010111101001000000", "0000000000100101001001100100101001000000", "0000000000100101001010010011100001001100", "0000000000111100001000100010001111000000", "0110010010100101001010010100100110000000", "0010001100001000010000100001000111000000", "0110010010000100010001000100001111000000", "0110010010000100110000010100100110000000", "0110010100101001010010100111100010000000", "1111010000100001110000010100100110000000", "0110010010100001110010010100100110000000", "1111000010000100010000100010000100000000", "0110010010100100110010010100100110000000", "0110010010100100111000010100100110000000", "0010000100001000010000100000000010000000", "0110010010000100010000100000000010000000", "0000000000000000000000000011000110000000", "0100000100000000110010010111101000001110", "0010001000000000110010010111101000001110", "0010000100010000000000000000000000000000", "0000010000110001110011110111001100010000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000", "0000000000000000000000000000000000000000");
  ATTRIBUTE RAM_STYLE : string;
  ATTRIBUTE RAM_STYLE of rom: signal is "BLOCK";

BEGIN

  PROCESS (CLOCK)
  BEGIN
    IF (CLOCK'event AND CLOCK = '1') THEN
      DATA_OUT <= STD_LOGIC_VECTOR( rom(to_integer(UNSIGNED(ADDR_R))) );
    END IF;
  END PROCESS;
  
END Behavioral;